  module forwarding (
  	input targetReg,
  	input targetData,
  	input MEM_reg,
  	input MEM_data,
  	input WB_reg,
  	input WB_data
  );
  
  endmodule