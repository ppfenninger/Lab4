module jumpTest (
	input[31:0] instruction,
	input[31:0] programCounter,
	output[31:0] jumpAddress,
	output doesJump
);

endmodule