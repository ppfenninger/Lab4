module jumpTest (
	input instruction,
	output jumpAddress,
	output doesJump
);

endmodule